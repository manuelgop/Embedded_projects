`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:52:42 02/10/2016 
// Design Name: 
// Module Name:    ProgCounter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ProgCounter(
    input PCIn,
    input Clk,
    input Cen,
    input Rst,
    output [7:0] PCOut
    );


endmodule
