`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:04:30 02/10/2016 
// Design Name: 
// Module Name:    Registers 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Registers(
    input [2:0] SelA,
    input [2:0] SelB,
    input [2:0] SelWR,
    input [7:0] Data,
    input Clk,
    input Cen,
    input Rst,
    input WE,
    output [7:0] OutA,
    output [7:0] OutB
    );


endmodule
