`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:01:01 02/10/2016 
// Design Name: 
// Module Name:    CtrlUnit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CtrlUnit(
    input [3:0] Oper,
    output [1:0] RegSrc_Op,
    output [2:0] ALUOp_Op,
    output RegWrite_Op,
    output Write7Seg_Op,
    output WriteLEDs_Op,
    output PCInc_Op,
    output Beq_Op,
    output [1:0] JiJr_Op
    );


endmodule
