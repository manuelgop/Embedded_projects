`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:10:52 02/10/2016 
// Design Name: 
// Module Name:    BrEq 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module BrEq(
    output M,
    input Sel,
    input InA,
    input InB
    );
	
	reg M;
	
	always@(*)
	begin 
		if (Sel)
			M = InB;
		else 
			M = InA;
	end
		
endmodule
